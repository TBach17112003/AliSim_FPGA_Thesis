library verilog;
use verilog.vl_types.all;
entity test_neoRNG is
end test_neoRNG;
