library verilog;
use verilog.vl_types.all;
entity test_RO is
end test_RO;
