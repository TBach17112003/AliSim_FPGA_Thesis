library verilog;
use verilog.vl_types.all;
entity test_Schedule is
end test_Schedule;
