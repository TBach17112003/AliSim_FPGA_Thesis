library verilog;
use verilog.vl_types.all;
entity PEran_tb is
end PEran_tb;
