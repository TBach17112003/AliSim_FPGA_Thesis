library verilog;
use verilog.vl_types.all;
entity moduleName is
end moduleName;
