library verilog;
use verilog.vl_types.all;
entity RG_tb is
end RG_tb;
