library verilog;
use verilog.vl_types.all;
entity PE_tb is
end PE_tb;
